module demux_1_2(
  input sel,
  input i,
  output y0,y1);
  assign y0=(~sel)&i;
  assign y1=sel&i;
endmodule
