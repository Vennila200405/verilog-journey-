module mux_4_1 (
  input  [1:0] sel,
  input  i0, i1, i2, i3,
  output y);
  assign y = sel[1] ? (sel[0] ? i3 : i2) :(sel[0] ? i1 : i0);
endmodule




















